library work;
use work.basicBuildingBlocksVhdl_package.all;